library IEEE;
use IEEE.STD_LOGIC_1164.ALL;	
use IEEE.NUMERIC_STD.ALL;
use WORK.lib_package.ALL;

entity datapath is
    port(
        rst, clk : in std_logic;
        K, N     : in unsigned(7 downto 0);

        -- counter control signals
        rst_i, inc_i : in std_logic;
        rst_j, inc_j : in std_logic;
        rst_m, inc_m : in std_logic;
        rst_n, inc_n : in std_logic;
        z_i, z_j, z_m, z_n : out std_logic;

        -- register controls
        rst_in, val_in_ld : in std_logic;
        rst_k, val_k_ld   : in std_logic;
        rst_sum, sum_ld   : in std_logic;


        -- memory signals
        base_in, base_k, base_out : in unsigned(17 downto 0);
        mem_addr_sel   : in std_logic_vector(1 downto 0);
        sum_sel        : in std_logic;
        mem_read_data  : in std_logic_vector(31 downto 0);
        mem_write_data : out std_logic_vector(31 downto 0);
        mem_addr       : out unsigned(17 downto 0)
    );
end datapath;

architecture rtl of datapath is
    -- signals
    signal S_sub_1, S, K_sub_1     : unsigned(7 downto 0):= (others => '0');
    signal i, j, m, n_out   : unsigned(7 downto 0) := (others => '0');
    signal val_in, val_k    : std_logic_vector(15 downto 0):= (others => '0');
    signal sum, sum_out, sum_in : std_logic_vector(31 downto 0):= (others => '0');
    signal addr_out, addr_in, addr_k : unsigned(17 downto 0):= (others => '0');

begin
    S       <= N - K + 1;

    -----------------------------------------------------------------
    -- COUNTERS
    -----------------------------------------------------------------
    i_up_counter : up_counter 
        
        port map (
            clk   => clk, 
            inc   => inc_i,
            rst   => rst_i,
            z     => z_i,
            count => i, 
            stop  => S
        );

    j_up_counter : up_counter 
        
        port map (
            clk   => clk, 
            inc   => inc_j,
            rst   => rst_j,
            z     => z_j,
            count => j, 
            stop  => S
        );

    m_up_counter : up_counter 
        
        port map (
            clk   => clk, 
            inc   => inc_m,
            rst   => rst_m,
            z     => z_m,
            count => m,
            stop  => K
        );

    n_up_counter : up_counter 
        
        port map (
            clk   => clk, 
            inc   => inc_n,
            rst   => rst_n,
            z     => z_n, 
            count => n_out,
            stop  => K
        );
    -----------------------------------------------------------------
    -- caculating address
    -----------------------------------------------------------------

addr_out <= base_out + resize(S * i + j, 18);
addr_in  <= base_in  + resize((j + n_out) + ((i + m) * N), 18);
addr_k   <= base_k   + resize((m * K) + n_out, 18);

mem_addr <= addr_out when mem_addr_sel = "00" else
            addr_in when mem_addr_sel = "01" else
            addr_k   when mem_addr_sel = "10" else
            (others => '0');


    -----------------------------------------------------------------
    -- REGISTERS
    -----------------------------------------------------------------
    val_in_reg : reg
        generic map ( DATA_WIDTH => 16 )
        port map (
            rst => rst_in,
            clk => clk,
            en  => val_in_ld,
            d   => mem_read_data(15 downto 0),
            q   => val_in
        );

    val_k_reg : reg
        generic map ( DATA_WIDTH => 16 )
        port map (
            rst => rst_k,
            clk => clk,
            en  => val_k_ld,
            d   => mem_read_data(15 downto 0),
            q   => val_k
        );

    sum_reg : reg
        generic map ( DATA_WIDTH => 32 )
        port map (
            rst => rst_sum,
            clk => clk,
            en  => sum_ld,
            d   => sum,
            q   => sum_out
        );

    -----------------------------------------------------------------
    -- calculating data
    -----------------------------------------------------------------
sum_in <= std_logic_vector(
    resize(signed(val_in) * signed(val_k), 32) + signed(sum_out)
);

    sum <= sum_in when sum_sel = '1' else (others => '0');
    mem_write_data <= sum_out;


end rtl;

